parameter coreConfig="RV32I";
parameter fetchWidth=4;
parameter GHRWidth=16;
parameter RASEntries=128;
parameter BTBEntries=4096;
parameter startPC='h00000000;
parameter FTQEntries=16;
parameter ROBEntries=64;
parameter architecturalRegCount=32;
parameter RATCheckpointCount=16;
parameter physicalRegCount=65;
parameter RSEntries=16;
parameter L1_instructionCacheWays=2;
parameter L1_instructionCacheSets=64;
parameter L1_instructionCacheBlockSizeBytes=32;
parameter ALUportCount=3;
parameter MEMportCount=1;
parameter FPUportCount=0;
parameter instruction_queue_depth=8;
parameter speculative=1;
parameter MOBEntries=16;
parameter dispatchWidth=4;
parameter commitWidth=4;
localparam physicalRegBits=$clog2(physicalRegCount);
localparam architecturalRegBits=$clog2(architecturalRegCount);
localparam RATCheckpointBits=$clog2(RATCheckpointCount);
