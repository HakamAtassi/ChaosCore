class dram_axi_agent extends cache_agent

    function new(string name, uvm_component parent);
        super.new(name, parent);
    endfunction

endclass