



module TL_magic_mem#(parameter bin = "";)(
    input logic clock,
    input logic reset,

    // Channel A


    // Channel D

);



endmodule