package instruction_cache_pkg;
    import uvm_pkg::*;


`include "cache_env.svh"
`include "cache_base_test.svh"

//agents
`include "cache_agent.svh"
`include "cpu_io_agent.svh"
`include "dram_axi_agent.svh"

`include "cache_req.svh"
`include "cpu_io_monitor.svh"
`include "cpu_io_driver.svh"


endpackage