parameter commitWidth=4;
parameter dispatchWidth=4;
parameter MOBEntries=16;
parameter speculative=true;
parameter instruction_queue_depth=8;
parameter FPUportCount=0;
parameter MEMportCount=1;
parameter ALUportCount=3;
parameter L1_instructionCacheBlockSizeBytes=32;
parameter L1_instructionCacheSets=64;
parameter L1_instructionCacheWays=2;
parameter RSEntries=16;
parameter physicalRegCount=65;
parameter RATCheckpointCount=16;
parameter architecturalRegCount=32;
parameter ROBEntries=64;
parameter FTQEntries=16;
parameter startPC="h00000000".U;
parameter BTBEntries=4096;
parameter RASEntries=128;
parameter GHRWidth=16;
parameter fetchWidth=4;
parameter coreConfig="RV32I";
