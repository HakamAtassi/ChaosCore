
module nReadmWrite (
      input  [5:0] raddr_0,
      input  [5:0] raddr_1,
      input  [5:0] raddr_2,
      input  [5:0] raddr_3,
      input  [5:0] raddr_4,
      input  [5:0] raddr_5,
      input  [5:0] raddr_6,
      input  [5:0] raddr_7,
      output [31:0] rdata_0,
      output [31:0] rdata_1,
      output [31:0] rdata_2,
      output [31:0] rdata_3,
      output [31:0] rdata_4,
      output [31:0] rdata_5,
      output [31:0] rdata_6,
      output [31:0] rdata_7,
      input  [5:0] waddr_0,
      input  [5:0] waddr_1,
      input  [5:0] waddr_2,
      input  [5:0] waddr_3,
      input   wen_0,
      input   wen_1,
      input   wen_2,
      input   wen_3,
      input  [31:0] wdata_0,
      input  [31:0] wdata_1,
      input  [31:0] wdata_2,
      input  [31:0] wdata_3,
      input   clock,
      input   reset);
  reg [31:0] _zz_72_;
  reg [31:0] _zz_73_;
  reg [31:0] _zz_74_;
  reg [31:0] _zz_75_;
  reg [31:0] _zz_76_;
  reg [31:0] _zz_77_;
  reg [31:0] _zz_78_;
  reg [31:0] _zz_79_;
  reg [31:0] _zz_80_;
  reg [31:0] _zz_81_;
  reg [31:0] _zz_82_;
  reg [31:0] _zz_83_;
  reg [31:0] _zz_84_;
  reg [31:0] _zz_85_;
  reg [31:0] _zz_86_;
  reg [31:0] _zz_87_;
  reg [31:0] _zz_88_;
  reg [31:0] _zz_89_;
  reg [31:0] _zz_90_;
  reg [31:0] _zz_91_;
  reg [31:0] _zz_92_;
  reg [31:0] _zz_93_;
  reg [31:0] _zz_94_;
  reg [31:0] _zz_95_;
  reg [31:0] _zz_96_;
  reg [31:0] _zz_97_;
  reg [31:0] _zz_98_;
  reg [31:0] _zz_99_;
  reg [31:0] _zz_100_;
  reg [31:0] _zz_101_;
  reg [31:0] _zz_102_;
  reg [31:0] _zz_103_;
  reg [1:0] _zz_104_;
  reg [1:0] _zz_105_;
  reg [1:0] _zz_106_;
  reg [1:0] _zz_107_;
  reg [1:0] _zz_108_;
  reg [1:0] _zz_109_;
  reg [1:0] _zz_110_;
  reg [1:0] _zz_111_;
  reg [31:0] _zz_112_;
  reg [31:0] _zz_113_;
  reg [31:0] _zz_114_;
  reg [31:0] _zz_115_;
  reg [31:0] _zz_116_;
  reg [31:0] _zz_117_;
  reg [31:0] _zz_118_;
  reg [31:0] _zz_119_;
  wire [5:0] _zz_120_;
  wire [5:0] _zz_121_;
  wire [5:0] _zz_122_;
  wire [5:0] _zz_123_;
  wire [5:0] _zz_124_;
  wire [5:0] _zz_125_;
  wire [5:0] _zz_126_;
  wire [5:0] _zz_127_;
  wire [0:0] _zz_128_;
  wire [1:0] _zz_129_;
  wire [1:0] _zz_130_;
  wire  _zz_131_;
  wire  _zz_132_;
  wire  _zz_133_;
  wire  _zz_134_;
  wire  _zz_135_;
  wire  _zz_136_;
  wire  _zz_137_;
  wire  _zz_138_;
  wire [31:0] _zz_139_;
  wire  _zz_140_;
  wire  _zz_141_;
  wire  _zz_142_;
  wire  _zz_143_;
  wire  _zz_144_;
  wire  _zz_145_;
  wire  _zz_146_;
  wire  _zz_147_;
  wire [31:0] _zz_148_;
  wire  _zz_149_;
  wire  _zz_150_;
  wire  _zz_151_;
  wire  _zz_152_;
  wire  _zz_153_;
  wire  _zz_154_;
  wire  _zz_155_;
  wire  _zz_156_;
  wire [31:0] _zz_157_;
  wire  _zz_158_;
  wire  _zz_159_;
  wire  _zz_160_;
  wire  _zz_161_;
  wire  _zz_162_;
  wire  _zz_163_;
  wire  _zz_164_;
  wire  _zz_165_;
  wire [31:0] _zz_166_;
  reg [1:0] _zz_1_;
  reg [1:0] _zz_2_;
  reg [1:0] _zz_3_;
  reg [1:0] _zz_4_;
  reg [1:0] _zz_5_;
  reg [1:0] _zz_6_;
  reg [1:0] _zz_7_;
  reg [1:0] _zz_8_;
  reg [1:0] _zz_9_;
  reg [1:0] _zz_10_;
  reg [1:0] _zz_11_;
  reg [1:0] _zz_12_;
  reg [1:0] _zz_13_;
  reg [1:0] _zz_14_;
  reg [1:0] _zz_15_;
  reg [1:0] _zz_16_;
  reg [1:0] _zz_17_;
  reg [1:0] _zz_18_;
  reg [1:0] _zz_19_;
  reg [1:0] _zz_20_;
  reg [1:0] _zz_21_;
  reg [1:0] _zz_22_;
  reg [1:0] _zz_23_;
  reg [1:0] _zz_24_;
  reg [1:0] _zz_25_;
  reg [1:0] _zz_26_;
  reg [1:0] _zz_27_;
  reg [1:0] _zz_28_;
  reg [1:0] _zz_29_;
  reg [1:0] _zz_30_;
  reg [1:0] _zz_31_;
  reg [1:0] _zz_32_;
  reg [1:0] _zz_33_;
  reg [1:0] _zz_34_;
  reg [1:0] _zz_35_;
  reg [1:0] _zz_36_;
  reg [1:0] _zz_37_;
  reg [1:0] _zz_38_;
  reg [1:0] _zz_39_;
  reg [1:0] _zz_40_;
  reg [1:0] _zz_41_;
  reg [1:0] _zz_42_;
  reg [1:0] _zz_43_;
  reg [1:0] _zz_44_;
  reg [1:0] _zz_45_;
  reg [1:0] _zz_46_;
  reg [1:0] _zz_47_;
  reg [1:0] _zz_48_;
  reg [1:0] _zz_49_;
  reg [1:0] _zz_50_;
  reg [1:0] _zz_51_;
  reg [1:0] _zz_52_;
  reg [1:0] _zz_53_;
  reg [1:0] _zz_54_;
  reg [1:0] _zz_55_;
  reg [1:0] _zz_56_;
  reg [1:0] _zz_57_;
  reg [1:0] _zz_58_;
  reg [1:0] _zz_59_;
  reg [1:0] _zz_60_;
  reg [1:0] _zz_61_;
  reg [1:0] _zz_62_;
  reg [1:0] _zz_63_;
  reg [1:0] _zz_64_;
  wire [31:0] reads_0_0;
  wire [31:0] reads_0_1;
  wire [31:0] reads_0_2;
  wire [31:0] reads_0_3;
  wire [31:0] reads_0_4;
  wire [31:0] reads_0_5;
  wire [31:0] reads_0_6;
  wire [31:0] reads_0_7;
  wire [31:0] reads_1_0;
  wire [31:0] reads_1_1;
  wire [31:0] reads_1_2;
  wire [31:0] reads_1_3;
  wire [31:0] reads_1_4;
  wire [31:0] reads_1_5;
  wire [31:0] reads_1_6;
  wire [31:0] reads_1_7;
  wire [31:0] reads_2_0;
  wire [31:0] reads_2_1;
  wire [31:0] reads_2_2;
  wire [31:0] reads_2_3;
  wire [31:0] reads_2_4;
  wire [31:0] reads_2_5;
  wire [31:0] reads_2_6;
  wire [31:0] reads_2_7;
  wire [31:0] reads_3_0;
  wire [31:0] reads_3_1;
  wire [31:0] reads_3_2;
  wire [31:0] reads_3_3;
  wire [31:0] reads_3_4;
  wire [31:0] reads_3_5;
  wire [31:0] reads_3_6;
  wire [31:0] reads_3_7;
  wire [1:0] lvr_0;
  wire [1:0] lvr_1;
  wire [1:0] lvr_2;
  wire [1:0] lvr_3;
  wire [1:0] lvr_4;
  wire [1:0] lvr_5;
  wire [1:0] lvr_6;
  wire [1:0] lvr_7;
  reg [1:0] banks_0;
  reg [1:0] banks_1;
  reg [1:0] banks_2;
  reg [1:0] banks_3;
  reg [1:0] banks_4;
  reg [1:0] banks_5;
  reg [1:0] banks_6;
  reg [1:0] banks_7;
  wire [63:0] _zz_65_;
  wire [63:0] _zz_66_;
  wire [1:0] _zz_67_;
  wire [63:0] _zz_68_;
  wire [1:0] _zz_69_;
  wire [63:0] _zz_70_;
  wire [1:0] _zz_71_;
  (* ramstyle = "no_rw_check, mlab" *) reg [31:0] rams_0 [0:63];
  (* ramstyle = "no_rw_check, mlab" *) reg [31:0] rams_1 [0:63];
  (* ramstyle = "no_rw_check, mlab" *) reg [31:0] rams_2 [0:63];
  (* ramstyle = "no_rw_check, mlab" *) reg [31:0] rams_3 [0:63];
  assign _zz_120_ = raddr_0;
  assign _zz_121_ = raddr_1;
  assign _zz_122_ = raddr_2;
  assign _zz_123_ = raddr_3;
  assign _zz_124_ = raddr_4;
  assign _zz_125_ = raddr_5;
  assign _zz_126_ = raddr_6;
  assign _zz_127_ = raddr_7;
  assign _zz_128_ = (1'b1);
  assign _zz_129_ = (2'b10);
  assign _zz_130_ = (2'b11);
  assign _zz_131_ = 1'b1;
  assign _zz_132_ = 1'b1;
  assign _zz_133_ = 1'b1;
  assign _zz_134_ = 1'b1;
  assign _zz_135_ = 1'b1;
  assign _zz_136_ = 1'b1;
  assign _zz_137_ = 1'b1;
  assign _zz_138_ = 1'b1;
  assign _zz_139_ = wdata_0;
  assign _zz_140_ = 1'b1;
  assign _zz_141_ = 1'b1;
  assign _zz_142_ = 1'b1;
  assign _zz_143_ = 1'b1;
  assign _zz_144_ = 1'b1;
  assign _zz_145_ = 1'b1;
  assign _zz_146_ = 1'b1;
  assign _zz_147_ = 1'b1;
  assign _zz_148_ = wdata_1;
  assign _zz_149_ = 1'b1;
  assign _zz_150_ = 1'b1;
  assign _zz_151_ = 1'b1;
  assign _zz_152_ = 1'b1;
  assign _zz_153_ = 1'b1;
  assign _zz_154_ = 1'b1;
  assign _zz_155_ = 1'b1;
  assign _zz_156_ = 1'b1;
  assign _zz_157_ = wdata_2;
  assign _zz_158_ = 1'b1;
  assign _zz_159_ = 1'b1;
  assign _zz_160_ = 1'b1;
  assign _zz_161_ = 1'b1;
  assign _zz_162_ = 1'b1;
  assign _zz_163_ = 1'b1;
  assign _zz_164_ = 1'b1;
  assign _zz_165_ = 1'b1;
  assign _zz_166_ = wdata_3;
  always @ (posedge clock) begin
    if(_zz_131_) begin
      _zz_72_ <= rams_0[raddr_0];
    end
  end

  always @ (posedge clock) begin
    if(_zz_132_) begin
      _zz_73_ <= rams_0[raddr_1];
    end
  end

  always @ (posedge clock) begin
    if(_zz_133_) begin
      _zz_74_ <= rams_0[raddr_2];
    end
  end

  always @ (posedge clock) begin
    if(_zz_134_) begin
      _zz_75_ <= rams_0[raddr_3];
    end
  end

  always @ (posedge clock) begin
    if(_zz_135_) begin
      _zz_76_ <= rams_0[raddr_4];
    end
  end

  always @ (posedge clock) begin
    if(_zz_136_) begin
      _zz_77_ <= rams_0[raddr_5];
    end
  end

  always @ (posedge clock) begin
    if(_zz_137_) begin
      _zz_78_ <= rams_0[raddr_6];
    end
  end

  always @ (posedge clock) begin
    if(_zz_138_) begin
      _zz_79_ <= rams_0[raddr_7];
    end
  end

  always @ (posedge clock) begin
    if(wen_0) begin
      rams_0[waddr_0] <= _zz_139_;
    end
  end

  always @ (posedge clock) begin
    if(_zz_140_) begin
      _zz_80_ <= rams_1[raddr_0];
    end
  end

  always @ (posedge clock) begin
    if(_zz_141_) begin
      _zz_81_ <= rams_1[raddr_1];
    end
  end

  always @ (posedge clock) begin
    if(_zz_142_) begin
      _zz_82_ <= rams_1[raddr_2];
    end
  end

  always @ (posedge clock) begin
    if(_zz_143_) begin
      _zz_83_ <= rams_1[raddr_3];
    end
  end

  always @ (posedge clock) begin
    if(_zz_144_) begin
      _zz_84_ <= rams_1[raddr_4];
    end
  end

  always @ (posedge clock) begin
    if(_zz_145_) begin
      _zz_85_ <= rams_1[raddr_5];
    end
  end

  always @ (posedge clock) begin
    if(_zz_146_) begin
      _zz_86_ <= rams_1[raddr_6];
    end
  end

  always @ (posedge clock) begin
    if(_zz_147_) begin
      _zz_87_ <= rams_1[raddr_7];
    end
  end

  always @ (posedge clock) begin
    if(wen_1) begin
      rams_1[waddr_1] <= _zz_148_;
    end
  end

  always @ (posedge clock) begin
    if(_zz_149_) begin
      _zz_88_ <= rams_2[raddr_0];
    end
  end

  always @ (posedge clock) begin
    if(_zz_150_) begin
      _zz_89_ <= rams_2[raddr_1];
    end
  end

  always @ (posedge clock) begin
    if(_zz_151_) begin
      _zz_90_ <= rams_2[raddr_2];
    end
  end

  always @ (posedge clock) begin
    if(_zz_152_) begin
      _zz_91_ <= rams_2[raddr_3];
    end
  end

  always @ (posedge clock) begin
    if(_zz_153_) begin
      _zz_92_ <= rams_2[raddr_4];
    end
  end

  always @ (posedge clock) begin
    if(_zz_154_) begin
      _zz_93_ <= rams_2[raddr_5];
    end
  end

  always @ (posedge clock) begin
    if(_zz_155_) begin
      _zz_94_ <= rams_2[raddr_6];
    end
  end

  always @ (posedge clock) begin
    if(_zz_156_) begin
      _zz_95_ <= rams_2[raddr_7];
    end
  end

  always @ (posedge clock) begin
    if(wen_2) begin
      rams_2[waddr_2] <= _zz_157_;
    end
  end

  always @ (posedge clock) begin
    if(_zz_158_) begin
      _zz_96_ <= rams_3[raddr_0];
    end
  end

  always @ (posedge clock) begin
    if(_zz_159_) begin
      _zz_97_ <= rams_3[raddr_1];
    end
  end

  always @ (posedge clock) begin
    if(_zz_160_) begin
      _zz_98_ <= rams_3[raddr_2];
    end
  end

  always @ (posedge clock) begin
    if(_zz_161_) begin
      _zz_99_ <= rams_3[raddr_3];
    end
  end

  always @ (posedge clock) begin
    if(_zz_162_) begin
      _zz_100_ <= rams_3[raddr_4];
    end
  end

  always @ (posedge clock) begin
    if(_zz_163_) begin
      _zz_101_ <= rams_3[raddr_5];
    end
  end

  always @ (posedge clock) begin
    if(_zz_164_) begin
      _zz_102_ <= rams_3[raddr_6];
    end
  end

  always @ (posedge clock) begin
    if(_zz_165_) begin
      _zz_103_ <= rams_3[raddr_7];
    end
  end

  always @ (posedge clock) begin
    if(wen_3) begin
      rams_3[waddr_3] <= _zz_166_;
    end
  end

  always @(*) begin
    case(_zz_120_)
      6'b000000 : begin
        _zz_104_ = _zz_1_;
      end
      6'b000001 : begin
        _zz_104_ = _zz_2_;
      end
      6'b000010 : begin
        _zz_104_ = _zz_3_;
      end
      6'b000011 : begin
        _zz_104_ = _zz_4_;
      end
      6'b000100 : begin
        _zz_104_ = _zz_5_;
      end
      6'b000101 : begin
        _zz_104_ = _zz_6_;
      end
      6'b000110 : begin
        _zz_104_ = _zz_7_;
      end
      6'b000111 : begin
        _zz_104_ = _zz_8_;
      end
      6'b001000 : begin
        _zz_104_ = _zz_9_;
      end
      6'b001001 : begin
        _zz_104_ = _zz_10_;
      end
      6'b001010 : begin
        _zz_104_ = _zz_11_;
      end
      6'b001011 : begin
        _zz_104_ = _zz_12_;
      end
      6'b001100 : begin
        _zz_104_ = _zz_13_;
      end
      6'b001101 : begin
        _zz_104_ = _zz_14_;
      end
      6'b001110 : begin
        _zz_104_ = _zz_15_;
      end
      6'b001111 : begin
        _zz_104_ = _zz_16_;
      end
      6'b010000 : begin
        _zz_104_ = _zz_17_;
      end
      6'b010001 : begin
        _zz_104_ = _zz_18_;
      end
      6'b010010 : begin
        _zz_104_ = _zz_19_;
      end
      6'b010011 : begin
        _zz_104_ = _zz_20_;
      end
      6'b010100 : begin
        _zz_104_ = _zz_21_;
      end
      6'b010101 : begin
        _zz_104_ = _zz_22_;
      end
      6'b010110 : begin
        _zz_104_ = _zz_23_;
      end
      6'b010111 : begin
        _zz_104_ = _zz_24_;
      end
      6'b011000 : begin
        _zz_104_ = _zz_25_;
      end
      6'b011001 : begin
        _zz_104_ = _zz_26_;
      end
      6'b011010 : begin
        _zz_104_ = _zz_27_;
      end
      6'b011011 : begin
        _zz_104_ = _zz_28_;
      end
      6'b011100 : begin
        _zz_104_ = _zz_29_;
      end
      6'b011101 : begin
        _zz_104_ = _zz_30_;
      end
      6'b011110 : begin
        _zz_104_ = _zz_31_;
      end
      6'b011111 : begin
        _zz_104_ = _zz_32_;
      end
      6'b100000 : begin
        _zz_104_ = _zz_33_;
      end
      6'b100001 : begin
        _zz_104_ = _zz_34_;
      end
      6'b100010 : begin
        _zz_104_ = _zz_35_;
      end
      6'b100011 : begin
        _zz_104_ = _zz_36_;
      end
      6'b100100 : begin
        _zz_104_ = _zz_37_;
      end
      6'b100101 : begin
        _zz_104_ = _zz_38_;
      end
      6'b100110 : begin
        _zz_104_ = _zz_39_;
      end
      6'b100111 : begin
        _zz_104_ = _zz_40_;
      end
      6'b101000 : begin
        _zz_104_ = _zz_41_;
      end
      6'b101001 : begin
        _zz_104_ = _zz_42_;
      end
      6'b101010 : begin
        _zz_104_ = _zz_43_;
      end
      6'b101011 : begin
        _zz_104_ = _zz_44_;
      end
      6'b101100 : begin
        _zz_104_ = _zz_45_;
      end
      6'b101101 : begin
        _zz_104_ = _zz_46_;
      end
      6'b101110 : begin
        _zz_104_ = _zz_47_;
      end
      6'b101111 : begin
        _zz_104_ = _zz_48_;
      end
      6'b110000 : begin
        _zz_104_ = _zz_49_;
      end
      6'b110001 : begin
        _zz_104_ = _zz_50_;
      end
      6'b110010 : begin
        _zz_104_ = _zz_51_;
      end
      6'b110011 : begin
        _zz_104_ = _zz_52_;
      end
      6'b110100 : begin
        _zz_104_ = _zz_53_;
      end
      6'b110101 : begin
        _zz_104_ = _zz_54_;
      end
      6'b110110 : begin
        _zz_104_ = _zz_55_;
      end
      6'b110111 : begin
        _zz_104_ = _zz_56_;
      end
      6'b111000 : begin
        _zz_104_ = _zz_57_;
      end
      6'b111001 : begin
        _zz_104_ = _zz_58_;
      end
      6'b111010 : begin
        _zz_104_ = _zz_59_;
      end
      6'b111011 : begin
        _zz_104_ = _zz_60_;
      end
      6'b111100 : begin
        _zz_104_ = _zz_61_;
      end
      6'b111101 : begin
        _zz_104_ = _zz_62_;
      end
      6'b111110 : begin
        _zz_104_ = _zz_63_;
      end
      default : begin
        _zz_104_ = _zz_64_;
      end
    endcase
  end

  always @(*) begin
    case(_zz_121_)
      6'b000000 : begin
        _zz_105_ = _zz_1_;
      end
      6'b000001 : begin
        _zz_105_ = _zz_2_;
      end
      6'b000010 : begin
        _zz_105_ = _zz_3_;
      end
      6'b000011 : begin
        _zz_105_ = _zz_4_;
      end
      6'b000100 : begin
        _zz_105_ = _zz_5_;
      end
      6'b000101 : begin
        _zz_105_ = _zz_6_;
      end
      6'b000110 : begin
        _zz_105_ = _zz_7_;
      end
      6'b000111 : begin
        _zz_105_ = _zz_8_;
      end
      6'b001000 : begin
        _zz_105_ = _zz_9_;
      end
      6'b001001 : begin
        _zz_105_ = _zz_10_;
      end
      6'b001010 : begin
        _zz_105_ = _zz_11_;
      end
      6'b001011 : begin
        _zz_105_ = _zz_12_;
      end
      6'b001100 : begin
        _zz_105_ = _zz_13_;
      end
      6'b001101 : begin
        _zz_105_ = _zz_14_;
      end
      6'b001110 : begin
        _zz_105_ = _zz_15_;
      end
      6'b001111 : begin
        _zz_105_ = _zz_16_;
      end
      6'b010000 : begin
        _zz_105_ = _zz_17_;
      end
      6'b010001 : begin
        _zz_105_ = _zz_18_;
      end
      6'b010010 : begin
        _zz_105_ = _zz_19_;
      end
      6'b010011 : begin
        _zz_105_ = _zz_20_;
      end
      6'b010100 : begin
        _zz_105_ = _zz_21_;
      end
      6'b010101 : begin
        _zz_105_ = _zz_22_;
      end
      6'b010110 : begin
        _zz_105_ = _zz_23_;
      end
      6'b010111 : begin
        _zz_105_ = _zz_24_;
      end
      6'b011000 : begin
        _zz_105_ = _zz_25_;
      end
      6'b011001 : begin
        _zz_105_ = _zz_26_;
      end
      6'b011010 : begin
        _zz_105_ = _zz_27_;
      end
      6'b011011 : begin
        _zz_105_ = _zz_28_;
      end
      6'b011100 : begin
        _zz_105_ = _zz_29_;
      end
      6'b011101 : begin
        _zz_105_ = _zz_30_;
      end
      6'b011110 : begin
        _zz_105_ = _zz_31_;
      end
      6'b011111 : begin
        _zz_105_ = _zz_32_;
      end
      6'b100000 : begin
        _zz_105_ = _zz_33_;
      end
      6'b100001 : begin
        _zz_105_ = _zz_34_;
      end
      6'b100010 : begin
        _zz_105_ = _zz_35_;
      end
      6'b100011 : begin
        _zz_105_ = _zz_36_;
      end
      6'b100100 : begin
        _zz_105_ = _zz_37_;
      end
      6'b100101 : begin
        _zz_105_ = _zz_38_;
      end
      6'b100110 : begin
        _zz_105_ = _zz_39_;
      end
      6'b100111 : begin
        _zz_105_ = _zz_40_;
      end
      6'b101000 : begin
        _zz_105_ = _zz_41_;
      end
      6'b101001 : begin
        _zz_105_ = _zz_42_;
      end
      6'b101010 : begin
        _zz_105_ = _zz_43_;
      end
      6'b101011 : begin
        _zz_105_ = _zz_44_;
      end
      6'b101100 : begin
        _zz_105_ = _zz_45_;
      end
      6'b101101 : begin
        _zz_105_ = _zz_46_;
      end
      6'b101110 : begin
        _zz_105_ = _zz_47_;
      end
      6'b101111 : begin
        _zz_105_ = _zz_48_;
      end
      6'b110000 : begin
        _zz_105_ = _zz_49_;
      end
      6'b110001 : begin
        _zz_105_ = _zz_50_;
      end
      6'b110010 : begin
        _zz_105_ = _zz_51_;
      end
      6'b110011 : begin
        _zz_105_ = _zz_52_;
      end
      6'b110100 : begin
        _zz_105_ = _zz_53_;
      end
      6'b110101 : begin
        _zz_105_ = _zz_54_;
      end
      6'b110110 : begin
        _zz_105_ = _zz_55_;
      end
      6'b110111 : begin
        _zz_105_ = _zz_56_;
      end
      6'b111000 : begin
        _zz_105_ = _zz_57_;
      end
      6'b111001 : begin
        _zz_105_ = _zz_58_;
      end
      6'b111010 : begin
        _zz_105_ = _zz_59_;
      end
      6'b111011 : begin
        _zz_105_ = _zz_60_;
      end
      6'b111100 : begin
        _zz_105_ = _zz_61_;
      end
      6'b111101 : begin
        _zz_105_ = _zz_62_;
      end
      6'b111110 : begin
        _zz_105_ = _zz_63_;
      end
      default : begin
        _zz_105_ = _zz_64_;
      end
    endcase
  end

  always @(*) begin
    case(_zz_122_)
      6'b000000 : begin
        _zz_106_ = _zz_1_;
      end
      6'b000001 : begin
        _zz_106_ = _zz_2_;
      end
      6'b000010 : begin
        _zz_106_ = _zz_3_;
      end
      6'b000011 : begin
        _zz_106_ = _zz_4_;
      end
      6'b000100 : begin
        _zz_106_ = _zz_5_;
      end
      6'b000101 : begin
        _zz_106_ = _zz_6_;
      end
      6'b000110 : begin
        _zz_106_ = _zz_7_;
      end
      6'b000111 : begin
        _zz_106_ = _zz_8_;
      end
      6'b001000 : begin
        _zz_106_ = _zz_9_;
      end
      6'b001001 : begin
        _zz_106_ = _zz_10_;
      end
      6'b001010 : begin
        _zz_106_ = _zz_11_;
      end
      6'b001011 : begin
        _zz_106_ = _zz_12_;
      end
      6'b001100 : begin
        _zz_106_ = _zz_13_;
      end
      6'b001101 : begin
        _zz_106_ = _zz_14_;
      end
      6'b001110 : begin
        _zz_106_ = _zz_15_;
      end
      6'b001111 : begin
        _zz_106_ = _zz_16_;
      end
      6'b010000 : begin
        _zz_106_ = _zz_17_;
      end
      6'b010001 : begin
        _zz_106_ = _zz_18_;
      end
      6'b010010 : begin
        _zz_106_ = _zz_19_;
      end
      6'b010011 : begin
        _zz_106_ = _zz_20_;
      end
      6'b010100 : begin
        _zz_106_ = _zz_21_;
      end
      6'b010101 : begin
        _zz_106_ = _zz_22_;
      end
      6'b010110 : begin
        _zz_106_ = _zz_23_;
      end
      6'b010111 : begin
        _zz_106_ = _zz_24_;
      end
      6'b011000 : begin
        _zz_106_ = _zz_25_;
      end
      6'b011001 : begin
        _zz_106_ = _zz_26_;
      end
      6'b011010 : begin
        _zz_106_ = _zz_27_;
      end
      6'b011011 : begin
        _zz_106_ = _zz_28_;
      end
      6'b011100 : begin
        _zz_106_ = _zz_29_;
      end
      6'b011101 : begin
        _zz_106_ = _zz_30_;
      end
      6'b011110 : begin
        _zz_106_ = _zz_31_;
      end
      6'b011111 : begin
        _zz_106_ = _zz_32_;
      end
      6'b100000 : begin
        _zz_106_ = _zz_33_;
      end
      6'b100001 : begin
        _zz_106_ = _zz_34_;
      end
      6'b100010 : begin
        _zz_106_ = _zz_35_;
      end
      6'b100011 : begin
        _zz_106_ = _zz_36_;
      end
      6'b100100 : begin
        _zz_106_ = _zz_37_;
      end
      6'b100101 : begin
        _zz_106_ = _zz_38_;
      end
      6'b100110 : begin
        _zz_106_ = _zz_39_;
      end
      6'b100111 : begin
        _zz_106_ = _zz_40_;
      end
      6'b101000 : begin
        _zz_106_ = _zz_41_;
      end
      6'b101001 : begin
        _zz_106_ = _zz_42_;
      end
      6'b101010 : begin
        _zz_106_ = _zz_43_;
      end
      6'b101011 : begin
        _zz_106_ = _zz_44_;
      end
      6'b101100 : begin
        _zz_106_ = _zz_45_;
      end
      6'b101101 : begin
        _zz_106_ = _zz_46_;
      end
      6'b101110 : begin
        _zz_106_ = _zz_47_;
      end
      6'b101111 : begin
        _zz_106_ = _zz_48_;
      end
      6'b110000 : begin
        _zz_106_ = _zz_49_;
      end
      6'b110001 : begin
        _zz_106_ = _zz_50_;
      end
      6'b110010 : begin
        _zz_106_ = _zz_51_;
      end
      6'b110011 : begin
        _zz_106_ = _zz_52_;
      end
      6'b110100 : begin
        _zz_106_ = _zz_53_;
      end
      6'b110101 : begin
        _zz_106_ = _zz_54_;
      end
      6'b110110 : begin
        _zz_106_ = _zz_55_;
      end
      6'b110111 : begin
        _zz_106_ = _zz_56_;
      end
      6'b111000 : begin
        _zz_106_ = _zz_57_;
      end
      6'b111001 : begin
        _zz_106_ = _zz_58_;
      end
      6'b111010 : begin
        _zz_106_ = _zz_59_;
      end
      6'b111011 : begin
        _zz_106_ = _zz_60_;
      end
      6'b111100 : begin
        _zz_106_ = _zz_61_;
      end
      6'b111101 : begin
        _zz_106_ = _zz_62_;
      end
      6'b111110 : begin
        _zz_106_ = _zz_63_;
      end
      default : begin
        _zz_106_ = _zz_64_;
      end
    endcase
  end

  always @(*) begin
    case(_zz_123_)
      6'b000000 : begin
        _zz_107_ = _zz_1_;
      end
      6'b000001 : begin
        _zz_107_ = _zz_2_;
      end
      6'b000010 : begin
        _zz_107_ = _zz_3_;
      end
      6'b000011 : begin
        _zz_107_ = _zz_4_;
      end
      6'b000100 : begin
        _zz_107_ = _zz_5_;
      end
      6'b000101 : begin
        _zz_107_ = _zz_6_;
      end
      6'b000110 : begin
        _zz_107_ = _zz_7_;
      end
      6'b000111 : begin
        _zz_107_ = _zz_8_;
      end
      6'b001000 : begin
        _zz_107_ = _zz_9_;
      end
      6'b001001 : begin
        _zz_107_ = _zz_10_;
      end
      6'b001010 : begin
        _zz_107_ = _zz_11_;
      end
      6'b001011 : begin
        _zz_107_ = _zz_12_;
      end
      6'b001100 : begin
        _zz_107_ = _zz_13_;
      end
      6'b001101 : begin
        _zz_107_ = _zz_14_;
      end
      6'b001110 : begin
        _zz_107_ = _zz_15_;
      end
      6'b001111 : begin
        _zz_107_ = _zz_16_;
      end
      6'b010000 : begin
        _zz_107_ = _zz_17_;
      end
      6'b010001 : begin
        _zz_107_ = _zz_18_;
      end
      6'b010010 : begin
        _zz_107_ = _zz_19_;
      end
      6'b010011 : begin
        _zz_107_ = _zz_20_;
      end
      6'b010100 : begin
        _zz_107_ = _zz_21_;
      end
      6'b010101 : begin
        _zz_107_ = _zz_22_;
      end
      6'b010110 : begin
        _zz_107_ = _zz_23_;
      end
      6'b010111 : begin
        _zz_107_ = _zz_24_;
      end
      6'b011000 : begin
        _zz_107_ = _zz_25_;
      end
      6'b011001 : begin
        _zz_107_ = _zz_26_;
      end
      6'b011010 : begin
        _zz_107_ = _zz_27_;
      end
      6'b011011 : begin
        _zz_107_ = _zz_28_;
      end
      6'b011100 : begin
        _zz_107_ = _zz_29_;
      end
      6'b011101 : begin
        _zz_107_ = _zz_30_;
      end
      6'b011110 : begin
        _zz_107_ = _zz_31_;
      end
      6'b011111 : begin
        _zz_107_ = _zz_32_;
      end
      6'b100000 : begin
        _zz_107_ = _zz_33_;
      end
      6'b100001 : begin
        _zz_107_ = _zz_34_;
      end
      6'b100010 : begin
        _zz_107_ = _zz_35_;
      end
      6'b100011 : begin
        _zz_107_ = _zz_36_;
      end
      6'b100100 : begin
        _zz_107_ = _zz_37_;
      end
      6'b100101 : begin
        _zz_107_ = _zz_38_;
      end
      6'b100110 : begin
        _zz_107_ = _zz_39_;
      end
      6'b100111 : begin
        _zz_107_ = _zz_40_;
      end
      6'b101000 : begin
        _zz_107_ = _zz_41_;
      end
      6'b101001 : begin
        _zz_107_ = _zz_42_;
      end
      6'b101010 : begin
        _zz_107_ = _zz_43_;
      end
      6'b101011 : begin
        _zz_107_ = _zz_44_;
      end
      6'b101100 : begin
        _zz_107_ = _zz_45_;
      end
      6'b101101 : begin
        _zz_107_ = _zz_46_;
      end
      6'b101110 : begin
        _zz_107_ = _zz_47_;
      end
      6'b101111 : begin
        _zz_107_ = _zz_48_;
      end
      6'b110000 : begin
        _zz_107_ = _zz_49_;
      end
      6'b110001 : begin
        _zz_107_ = _zz_50_;
      end
      6'b110010 : begin
        _zz_107_ = _zz_51_;
      end
      6'b110011 : begin
        _zz_107_ = _zz_52_;
      end
      6'b110100 : begin
        _zz_107_ = _zz_53_;
      end
      6'b110101 : begin
        _zz_107_ = _zz_54_;
      end
      6'b110110 : begin
        _zz_107_ = _zz_55_;
      end
      6'b110111 : begin
        _zz_107_ = _zz_56_;
      end
      6'b111000 : begin
        _zz_107_ = _zz_57_;
      end
      6'b111001 : begin
        _zz_107_ = _zz_58_;
      end
      6'b111010 : begin
        _zz_107_ = _zz_59_;
      end
      6'b111011 : begin
        _zz_107_ = _zz_60_;
      end
      6'b111100 : begin
        _zz_107_ = _zz_61_;
      end
      6'b111101 : begin
        _zz_107_ = _zz_62_;
      end
      6'b111110 : begin
        _zz_107_ = _zz_63_;
      end
      default : begin
        _zz_107_ = _zz_64_;
      end
    endcase
  end

  always @(*) begin
    case(_zz_124_)
      6'b000000 : begin
        _zz_108_ = _zz_1_;
      end
      6'b000001 : begin
        _zz_108_ = _zz_2_;
      end
      6'b000010 : begin
        _zz_108_ = _zz_3_;
      end
      6'b000011 : begin
        _zz_108_ = _zz_4_;
      end
      6'b000100 : begin
        _zz_108_ = _zz_5_;
      end
      6'b000101 : begin
        _zz_108_ = _zz_6_;
      end
      6'b000110 : begin
        _zz_108_ = _zz_7_;
      end
      6'b000111 : begin
        _zz_108_ = _zz_8_;
      end
      6'b001000 : begin
        _zz_108_ = _zz_9_;
      end
      6'b001001 : begin
        _zz_108_ = _zz_10_;
      end
      6'b001010 : begin
        _zz_108_ = _zz_11_;
      end
      6'b001011 : begin
        _zz_108_ = _zz_12_;
      end
      6'b001100 : begin
        _zz_108_ = _zz_13_;
      end
      6'b001101 : begin
        _zz_108_ = _zz_14_;
      end
      6'b001110 : begin
        _zz_108_ = _zz_15_;
      end
      6'b001111 : begin
        _zz_108_ = _zz_16_;
      end
      6'b010000 : begin
        _zz_108_ = _zz_17_;
      end
      6'b010001 : begin
        _zz_108_ = _zz_18_;
      end
      6'b010010 : begin
        _zz_108_ = _zz_19_;
      end
      6'b010011 : begin
        _zz_108_ = _zz_20_;
      end
      6'b010100 : begin
        _zz_108_ = _zz_21_;
      end
      6'b010101 : begin
        _zz_108_ = _zz_22_;
      end
      6'b010110 : begin
        _zz_108_ = _zz_23_;
      end
      6'b010111 : begin
        _zz_108_ = _zz_24_;
      end
      6'b011000 : begin
        _zz_108_ = _zz_25_;
      end
      6'b011001 : begin
        _zz_108_ = _zz_26_;
      end
      6'b011010 : begin
        _zz_108_ = _zz_27_;
      end
      6'b011011 : begin
        _zz_108_ = _zz_28_;
      end
      6'b011100 : begin
        _zz_108_ = _zz_29_;
      end
      6'b011101 : begin
        _zz_108_ = _zz_30_;
      end
      6'b011110 : begin
        _zz_108_ = _zz_31_;
      end
      6'b011111 : begin
        _zz_108_ = _zz_32_;
      end
      6'b100000 : begin
        _zz_108_ = _zz_33_;
      end
      6'b100001 : begin
        _zz_108_ = _zz_34_;
      end
      6'b100010 : begin
        _zz_108_ = _zz_35_;
      end
      6'b100011 : begin
        _zz_108_ = _zz_36_;
      end
      6'b100100 : begin
        _zz_108_ = _zz_37_;
      end
      6'b100101 : begin
        _zz_108_ = _zz_38_;
      end
      6'b100110 : begin
        _zz_108_ = _zz_39_;
      end
      6'b100111 : begin
        _zz_108_ = _zz_40_;
      end
      6'b101000 : begin
        _zz_108_ = _zz_41_;
      end
      6'b101001 : begin
        _zz_108_ = _zz_42_;
      end
      6'b101010 : begin
        _zz_108_ = _zz_43_;
      end
      6'b101011 : begin
        _zz_108_ = _zz_44_;
      end
      6'b101100 : begin
        _zz_108_ = _zz_45_;
      end
      6'b101101 : begin
        _zz_108_ = _zz_46_;
      end
      6'b101110 : begin
        _zz_108_ = _zz_47_;
      end
      6'b101111 : begin
        _zz_108_ = _zz_48_;
      end
      6'b110000 : begin
        _zz_108_ = _zz_49_;
      end
      6'b110001 : begin
        _zz_108_ = _zz_50_;
      end
      6'b110010 : begin
        _zz_108_ = _zz_51_;
      end
      6'b110011 : begin
        _zz_108_ = _zz_52_;
      end
      6'b110100 : begin
        _zz_108_ = _zz_53_;
      end
      6'b110101 : begin
        _zz_108_ = _zz_54_;
      end
      6'b110110 : begin
        _zz_108_ = _zz_55_;
      end
      6'b110111 : begin
        _zz_108_ = _zz_56_;
      end
      6'b111000 : begin
        _zz_108_ = _zz_57_;
      end
      6'b111001 : begin
        _zz_108_ = _zz_58_;
      end
      6'b111010 : begin
        _zz_108_ = _zz_59_;
      end
      6'b111011 : begin
        _zz_108_ = _zz_60_;
      end
      6'b111100 : begin
        _zz_108_ = _zz_61_;
      end
      6'b111101 : begin
        _zz_108_ = _zz_62_;
      end
      6'b111110 : begin
        _zz_108_ = _zz_63_;
      end
      default : begin
        _zz_108_ = _zz_64_;
      end
    endcase
  end

  always @(*) begin
    case(_zz_125_)
      6'b000000 : begin
        _zz_109_ = _zz_1_;
      end
      6'b000001 : begin
        _zz_109_ = _zz_2_;
      end
      6'b000010 : begin
        _zz_109_ = _zz_3_;
      end
      6'b000011 : begin
        _zz_109_ = _zz_4_;
      end
      6'b000100 : begin
        _zz_109_ = _zz_5_;
      end
      6'b000101 : begin
        _zz_109_ = _zz_6_;
      end
      6'b000110 : begin
        _zz_109_ = _zz_7_;
      end
      6'b000111 : begin
        _zz_109_ = _zz_8_;
      end
      6'b001000 : begin
        _zz_109_ = _zz_9_;
      end
      6'b001001 : begin
        _zz_109_ = _zz_10_;
      end
      6'b001010 : begin
        _zz_109_ = _zz_11_;
      end
      6'b001011 : begin
        _zz_109_ = _zz_12_;
      end
      6'b001100 : begin
        _zz_109_ = _zz_13_;
      end
      6'b001101 : begin
        _zz_109_ = _zz_14_;
      end
      6'b001110 : begin
        _zz_109_ = _zz_15_;
      end
      6'b001111 : begin
        _zz_109_ = _zz_16_;
      end
      6'b010000 : begin
        _zz_109_ = _zz_17_;
      end
      6'b010001 : begin
        _zz_109_ = _zz_18_;
      end
      6'b010010 : begin
        _zz_109_ = _zz_19_;
      end
      6'b010011 : begin
        _zz_109_ = _zz_20_;
      end
      6'b010100 : begin
        _zz_109_ = _zz_21_;
      end
      6'b010101 : begin
        _zz_109_ = _zz_22_;
      end
      6'b010110 : begin
        _zz_109_ = _zz_23_;
      end
      6'b010111 : begin
        _zz_109_ = _zz_24_;
      end
      6'b011000 : begin
        _zz_109_ = _zz_25_;
      end
      6'b011001 : begin
        _zz_109_ = _zz_26_;
      end
      6'b011010 : begin
        _zz_109_ = _zz_27_;
      end
      6'b011011 : begin
        _zz_109_ = _zz_28_;
      end
      6'b011100 : begin
        _zz_109_ = _zz_29_;
      end
      6'b011101 : begin
        _zz_109_ = _zz_30_;
      end
      6'b011110 : begin
        _zz_109_ = _zz_31_;
      end
      6'b011111 : begin
        _zz_109_ = _zz_32_;
      end
      6'b100000 : begin
        _zz_109_ = _zz_33_;
      end
      6'b100001 : begin
        _zz_109_ = _zz_34_;
      end
      6'b100010 : begin
        _zz_109_ = _zz_35_;
      end
      6'b100011 : begin
        _zz_109_ = _zz_36_;
      end
      6'b100100 : begin
        _zz_109_ = _zz_37_;
      end
      6'b100101 : begin
        _zz_109_ = _zz_38_;
      end
      6'b100110 : begin
        _zz_109_ = _zz_39_;
      end
      6'b100111 : begin
        _zz_109_ = _zz_40_;
      end
      6'b101000 : begin
        _zz_109_ = _zz_41_;
      end
      6'b101001 : begin
        _zz_109_ = _zz_42_;
      end
      6'b101010 : begin
        _zz_109_ = _zz_43_;
      end
      6'b101011 : begin
        _zz_109_ = _zz_44_;
      end
      6'b101100 : begin
        _zz_109_ = _zz_45_;
      end
      6'b101101 : begin
        _zz_109_ = _zz_46_;
      end
      6'b101110 : begin
        _zz_109_ = _zz_47_;
      end
      6'b101111 : begin
        _zz_109_ = _zz_48_;
      end
      6'b110000 : begin
        _zz_109_ = _zz_49_;
      end
      6'b110001 : begin
        _zz_109_ = _zz_50_;
      end
      6'b110010 : begin
        _zz_109_ = _zz_51_;
      end
      6'b110011 : begin
        _zz_109_ = _zz_52_;
      end
      6'b110100 : begin
        _zz_109_ = _zz_53_;
      end
      6'b110101 : begin
        _zz_109_ = _zz_54_;
      end
      6'b110110 : begin
        _zz_109_ = _zz_55_;
      end
      6'b110111 : begin
        _zz_109_ = _zz_56_;
      end
      6'b111000 : begin
        _zz_109_ = _zz_57_;
      end
      6'b111001 : begin
        _zz_109_ = _zz_58_;
      end
      6'b111010 : begin
        _zz_109_ = _zz_59_;
      end
      6'b111011 : begin
        _zz_109_ = _zz_60_;
      end
      6'b111100 : begin
        _zz_109_ = _zz_61_;
      end
      6'b111101 : begin
        _zz_109_ = _zz_62_;
      end
      6'b111110 : begin
        _zz_109_ = _zz_63_;
      end
      default : begin
        _zz_109_ = _zz_64_;
      end
    endcase
  end

  always @(*) begin
    case(_zz_126_)
      6'b000000 : begin
        _zz_110_ = _zz_1_;
      end
      6'b000001 : begin
        _zz_110_ = _zz_2_;
      end
      6'b000010 : begin
        _zz_110_ = _zz_3_;
      end
      6'b000011 : begin
        _zz_110_ = _zz_4_;
      end
      6'b000100 : begin
        _zz_110_ = _zz_5_;
      end
      6'b000101 : begin
        _zz_110_ = _zz_6_;
      end
      6'b000110 : begin
        _zz_110_ = _zz_7_;
      end
      6'b000111 : begin
        _zz_110_ = _zz_8_;
      end
      6'b001000 : begin
        _zz_110_ = _zz_9_;
      end
      6'b001001 : begin
        _zz_110_ = _zz_10_;
      end
      6'b001010 : begin
        _zz_110_ = _zz_11_;
      end
      6'b001011 : begin
        _zz_110_ = _zz_12_;
      end
      6'b001100 : begin
        _zz_110_ = _zz_13_;
      end
      6'b001101 : begin
        _zz_110_ = _zz_14_;
      end
      6'b001110 : begin
        _zz_110_ = _zz_15_;
      end
      6'b001111 : begin
        _zz_110_ = _zz_16_;
      end
      6'b010000 : begin
        _zz_110_ = _zz_17_;
      end
      6'b010001 : begin
        _zz_110_ = _zz_18_;
      end
      6'b010010 : begin
        _zz_110_ = _zz_19_;
      end
      6'b010011 : begin
        _zz_110_ = _zz_20_;
      end
      6'b010100 : begin
        _zz_110_ = _zz_21_;
      end
      6'b010101 : begin
        _zz_110_ = _zz_22_;
      end
      6'b010110 : begin
        _zz_110_ = _zz_23_;
      end
      6'b010111 : begin
        _zz_110_ = _zz_24_;
      end
      6'b011000 : begin
        _zz_110_ = _zz_25_;
      end
      6'b011001 : begin
        _zz_110_ = _zz_26_;
      end
      6'b011010 : begin
        _zz_110_ = _zz_27_;
      end
      6'b011011 : begin
        _zz_110_ = _zz_28_;
      end
      6'b011100 : begin
        _zz_110_ = _zz_29_;
      end
      6'b011101 : begin
        _zz_110_ = _zz_30_;
      end
      6'b011110 : begin
        _zz_110_ = _zz_31_;
      end
      6'b011111 : begin
        _zz_110_ = _zz_32_;
      end
      6'b100000 : begin
        _zz_110_ = _zz_33_;
      end
      6'b100001 : begin
        _zz_110_ = _zz_34_;
      end
      6'b100010 : begin
        _zz_110_ = _zz_35_;
      end
      6'b100011 : begin
        _zz_110_ = _zz_36_;
      end
      6'b100100 : begin
        _zz_110_ = _zz_37_;
      end
      6'b100101 : begin
        _zz_110_ = _zz_38_;
      end
      6'b100110 : begin
        _zz_110_ = _zz_39_;
      end
      6'b100111 : begin
        _zz_110_ = _zz_40_;
      end
      6'b101000 : begin
        _zz_110_ = _zz_41_;
      end
      6'b101001 : begin
        _zz_110_ = _zz_42_;
      end
      6'b101010 : begin
        _zz_110_ = _zz_43_;
      end
      6'b101011 : begin
        _zz_110_ = _zz_44_;
      end
      6'b101100 : begin
        _zz_110_ = _zz_45_;
      end
      6'b101101 : begin
        _zz_110_ = _zz_46_;
      end
      6'b101110 : begin
        _zz_110_ = _zz_47_;
      end
      6'b101111 : begin
        _zz_110_ = _zz_48_;
      end
      6'b110000 : begin
        _zz_110_ = _zz_49_;
      end
      6'b110001 : begin
        _zz_110_ = _zz_50_;
      end
      6'b110010 : begin
        _zz_110_ = _zz_51_;
      end
      6'b110011 : begin
        _zz_110_ = _zz_52_;
      end
      6'b110100 : begin
        _zz_110_ = _zz_53_;
      end
      6'b110101 : begin
        _zz_110_ = _zz_54_;
      end
      6'b110110 : begin
        _zz_110_ = _zz_55_;
      end
      6'b110111 : begin
        _zz_110_ = _zz_56_;
      end
      6'b111000 : begin
        _zz_110_ = _zz_57_;
      end
      6'b111001 : begin
        _zz_110_ = _zz_58_;
      end
      6'b111010 : begin
        _zz_110_ = _zz_59_;
      end
      6'b111011 : begin
        _zz_110_ = _zz_60_;
      end
      6'b111100 : begin
        _zz_110_ = _zz_61_;
      end
      6'b111101 : begin
        _zz_110_ = _zz_62_;
      end
      6'b111110 : begin
        _zz_110_ = _zz_63_;
      end
      default : begin
        _zz_110_ = _zz_64_;
      end
    endcase
  end

  always @(*) begin
    case(_zz_127_)
      6'b000000 : begin
        _zz_111_ = _zz_1_;
      end
      6'b000001 : begin
        _zz_111_ = _zz_2_;
      end
      6'b000010 : begin
        _zz_111_ = _zz_3_;
      end
      6'b000011 : begin
        _zz_111_ = _zz_4_;
      end
      6'b000100 : begin
        _zz_111_ = _zz_5_;
      end
      6'b000101 : begin
        _zz_111_ = _zz_6_;
      end
      6'b000110 : begin
        _zz_111_ = _zz_7_;
      end
      6'b000111 : begin
        _zz_111_ = _zz_8_;
      end
      6'b001000 : begin
        _zz_111_ = _zz_9_;
      end
      6'b001001 : begin
        _zz_111_ = _zz_10_;
      end
      6'b001010 : begin
        _zz_111_ = _zz_11_;
      end
      6'b001011 : begin
        _zz_111_ = _zz_12_;
      end
      6'b001100 : begin
        _zz_111_ = _zz_13_;
      end
      6'b001101 : begin
        _zz_111_ = _zz_14_;
      end
      6'b001110 : begin
        _zz_111_ = _zz_15_;
      end
      6'b001111 : begin
        _zz_111_ = _zz_16_;
      end
      6'b010000 : begin
        _zz_111_ = _zz_17_;
      end
      6'b010001 : begin
        _zz_111_ = _zz_18_;
      end
      6'b010010 : begin
        _zz_111_ = _zz_19_;
      end
      6'b010011 : begin
        _zz_111_ = _zz_20_;
      end
      6'b010100 : begin
        _zz_111_ = _zz_21_;
      end
      6'b010101 : begin
        _zz_111_ = _zz_22_;
      end
      6'b010110 : begin
        _zz_111_ = _zz_23_;
      end
      6'b010111 : begin
        _zz_111_ = _zz_24_;
      end
      6'b011000 : begin
        _zz_111_ = _zz_25_;
      end
      6'b011001 : begin
        _zz_111_ = _zz_26_;
      end
      6'b011010 : begin
        _zz_111_ = _zz_27_;
      end
      6'b011011 : begin
        _zz_111_ = _zz_28_;
      end
      6'b011100 : begin
        _zz_111_ = _zz_29_;
      end
      6'b011101 : begin
        _zz_111_ = _zz_30_;
      end
      6'b011110 : begin
        _zz_111_ = _zz_31_;
      end
      6'b011111 : begin
        _zz_111_ = _zz_32_;
      end
      6'b100000 : begin
        _zz_111_ = _zz_33_;
      end
      6'b100001 : begin
        _zz_111_ = _zz_34_;
      end
      6'b100010 : begin
        _zz_111_ = _zz_35_;
      end
      6'b100011 : begin
        _zz_111_ = _zz_36_;
      end
      6'b100100 : begin
        _zz_111_ = _zz_37_;
      end
      6'b100101 : begin
        _zz_111_ = _zz_38_;
      end
      6'b100110 : begin
        _zz_111_ = _zz_39_;
      end
      6'b100111 : begin
        _zz_111_ = _zz_40_;
      end
      6'b101000 : begin
        _zz_111_ = _zz_41_;
      end
      6'b101001 : begin
        _zz_111_ = _zz_42_;
      end
      6'b101010 : begin
        _zz_111_ = _zz_43_;
      end
      6'b101011 : begin
        _zz_111_ = _zz_44_;
      end
      6'b101100 : begin
        _zz_111_ = _zz_45_;
      end
      6'b101101 : begin
        _zz_111_ = _zz_46_;
      end
      6'b101110 : begin
        _zz_111_ = _zz_47_;
      end
      6'b101111 : begin
        _zz_111_ = _zz_48_;
      end
      6'b110000 : begin
        _zz_111_ = _zz_49_;
      end
      6'b110001 : begin
        _zz_111_ = _zz_50_;
      end
      6'b110010 : begin
        _zz_111_ = _zz_51_;
      end
      6'b110011 : begin
        _zz_111_ = _zz_52_;
      end
      6'b110100 : begin
        _zz_111_ = _zz_53_;
      end
      6'b110101 : begin
        _zz_111_ = _zz_54_;
      end
      6'b110110 : begin
        _zz_111_ = _zz_55_;
      end
      6'b110111 : begin
        _zz_111_ = _zz_56_;
      end
      6'b111000 : begin
        _zz_111_ = _zz_57_;
      end
      6'b111001 : begin
        _zz_111_ = _zz_58_;
      end
      6'b111010 : begin
        _zz_111_ = _zz_59_;
      end
      6'b111011 : begin
        _zz_111_ = _zz_60_;
      end
      6'b111100 : begin
        _zz_111_ = _zz_61_;
      end
      6'b111101 : begin
        _zz_111_ = _zz_62_;
      end
      6'b111110 : begin
        _zz_111_ = _zz_63_;
      end
      default : begin
        _zz_111_ = _zz_64_;
      end
    endcase
  end

  always @(*) begin
    case(banks_0)
      2'b00 : begin
        _zz_112_ = reads_0_0;
      end
      2'b01 : begin
        _zz_112_ = reads_1_0;
      end
      2'b10 : begin
        _zz_112_ = reads_2_0;
      end
      default : begin
        _zz_112_ = reads_3_0;
      end
    endcase
  end

  always @(*) begin
    case(banks_1)
      2'b00 : begin
        _zz_113_ = reads_0_1;
      end
      2'b01 : begin
        _zz_113_ = reads_1_1;
      end
      2'b10 : begin
        _zz_113_ = reads_2_1;
      end
      default : begin
        _zz_113_ = reads_3_1;
      end
    endcase
  end

  always @(*) begin
    case(banks_2)
      2'b00 : begin
        _zz_114_ = reads_0_2;
      end
      2'b01 : begin
        _zz_114_ = reads_1_2;
      end
      2'b10 : begin
        _zz_114_ = reads_2_2;
      end
      default : begin
        _zz_114_ = reads_3_2;
      end
    endcase
  end

  always @(*) begin
    case(banks_3)
      2'b00 : begin
        _zz_115_ = reads_0_3;
      end
      2'b01 : begin
        _zz_115_ = reads_1_3;
      end
      2'b10 : begin
        _zz_115_ = reads_2_3;
      end
      default : begin
        _zz_115_ = reads_3_3;
      end
    endcase
  end

  always @(*) begin
    case(banks_4)
      2'b00 : begin
        _zz_116_ = reads_0_4;
      end
      2'b01 : begin
        _zz_116_ = reads_1_4;
      end
      2'b10 : begin
        _zz_116_ = reads_2_4;
      end
      default : begin
        _zz_116_ = reads_3_4;
      end
    endcase
  end

  always @(*) begin
    case(banks_5)
      2'b00 : begin
        _zz_117_ = reads_0_5;
      end
      2'b01 : begin
        _zz_117_ = reads_1_5;
      end
      2'b10 : begin
        _zz_117_ = reads_2_5;
      end
      default : begin
        _zz_117_ = reads_3_5;
      end
    endcase
  end

  always @(*) begin
    case(banks_6)
      2'b00 : begin
        _zz_118_ = reads_0_6;
      end
      2'b01 : begin
        _zz_118_ = reads_1_6;
      end
      2'b10 : begin
        _zz_118_ = reads_2_6;
      end
      default : begin
        _zz_118_ = reads_3_6;
      end
    endcase
  end

  always @(*) begin
    case(banks_7)
      2'b00 : begin
        _zz_119_ = reads_0_7;
      end
      2'b01 : begin
        _zz_119_ = reads_1_7;
      end
      2'b10 : begin
        _zz_119_ = reads_2_7;
      end
      default : begin
        _zz_119_ = reads_3_7;
      end
    endcase
  end

  assign reads_0_0 = _zz_72_;
  assign reads_0_1 = _zz_73_;
  assign reads_0_2 = _zz_74_;
  assign reads_0_3 = _zz_75_;
  assign reads_0_4 = _zz_76_;
  assign reads_0_5 = _zz_77_;
  assign reads_0_6 = _zz_78_;
  assign reads_0_7 = _zz_79_;
  assign reads_1_0 = _zz_80_;
  assign reads_1_1 = _zz_81_;
  assign reads_1_2 = _zz_82_;
  assign reads_1_3 = _zz_83_;
  assign reads_1_4 = _zz_84_;
  assign reads_1_5 = _zz_85_;
  assign reads_1_6 = _zz_86_;
  assign reads_1_7 = _zz_87_;
  assign reads_2_0 = _zz_88_;
  assign reads_2_1 = _zz_89_;
  assign reads_2_2 = _zz_90_;
  assign reads_2_3 = _zz_91_;
  assign reads_2_4 = _zz_92_;
  assign reads_2_5 = _zz_93_;
  assign reads_2_6 = _zz_94_;
  assign reads_2_7 = _zz_95_;
  assign reads_3_0 = _zz_96_;
  assign reads_3_1 = _zz_97_;
  assign reads_3_2 = _zz_98_;
  assign reads_3_3 = _zz_99_;
  assign reads_3_4 = _zz_100_;
  assign reads_3_5 = _zz_101_;
  assign reads_3_6 = _zz_102_;
  assign reads_3_7 = _zz_103_;
  assign lvr_0 = _zz_104_;
  assign lvr_1 = _zz_105_;
  assign lvr_2 = _zz_106_;
  assign lvr_3 = _zz_107_;
  assign lvr_4 = _zz_108_;
  assign lvr_5 = _zz_109_;
  assign lvr_6 = _zz_110_;
  assign lvr_7 = _zz_111_;
  assign rdata_0 = _zz_112_;
  assign rdata_1 = _zz_113_;
  assign rdata_2 = _zz_114_;
  assign rdata_3 = _zz_115_;
  assign rdata_4 = _zz_116_;
  assign rdata_5 = _zz_117_;
  assign rdata_6 = _zz_118_;
  assign rdata_7 = _zz_119_;
  assign _zz_65_ = ({63'd0,(1'b1)} <<< waddr_0);
  assign _zz_66_ = ({63'd0,(1'b1)} <<< waddr_1);
  assign _zz_67_ = {1'd0, _zz_128_};
  assign _zz_68_ = ({63'd0,(1'b1)} <<< waddr_2);
  assign _zz_69_ = _zz_129_;
  assign _zz_70_ = ({63'd0,(1'b1)} <<< waddr_3);
  assign _zz_71_ = _zz_130_;
  always @ (posedge clock) begin
    banks_0 <= lvr_0;
    banks_1 <= lvr_1;
    banks_2 <= lvr_2;
    banks_3 <= lvr_3;
    banks_4 <= lvr_4;
    banks_5 <= lvr_5;
    banks_6 <= lvr_6;
    banks_7 <= lvr_7;
    if(wen_0)begin
      if(_zz_65_[0])begin
        _zz_1_ <= (2'b00);
      end
      if(_zz_65_[1])begin
        _zz_2_ <= (2'b00);
      end
      if(_zz_65_[2])begin
        _zz_3_ <= (2'b00);
      end
      if(_zz_65_[3])begin
        _zz_4_ <= (2'b00);
      end
      if(_zz_65_[4])begin
        _zz_5_ <= (2'b00);
      end
      if(_zz_65_[5])begin
        _zz_6_ <= (2'b00);
      end
      if(_zz_65_[6])begin
        _zz_7_ <= (2'b00);
      end
      if(_zz_65_[7])begin
        _zz_8_ <= (2'b00);
      end
      if(_zz_65_[8])begin
        _zz_9_ <= (2'b00);
      end
      if(_zz_65_[9])begin
        _zz_10_ <= (2'b00);
      end
      if(_zz_65_[10])begin
        _zz_11_ <= (2'b00);
      end
      if(_zz_65_[11])begin
        _zz_12_ <= (2'b00);
      end
      if(_zz_65_[12])begin
        _zz_13_ <= (2'b00);
      end
      if(_zz_65_[13])begin
        _zz_14_ <= (2'b00);
      end
      if(_zz_65_[14])begin
        _zz_15_ <= (2'b00);
      end
      if(_zz_65_[15])begin
        _zz_16_ <= (2'b00);
      end
      if(_zz_65_[16])begin
        _zz_17_ <= (2'b00);
      end
      if(_zz_65_[17])begin
        _zz_18_ <= (2'b00);
      end
      if(_zz_65_[18])begin
        _zz_19_ <= (2'b00);
      end
      if(_zz_65_[19])begin
        _zz_20_ <= (2'b00);
      end
      if(_zz_65_[20])begin
        _zz_21_ <= (2'b00);
      end
      if(_zz_65_[21])begin
        _zz_22_ <= (2'b00);
      end
      if(_zz_65_[22])begin
        _zz_23_ <= (2'b00);
      end
      if(_zz_65_[23])begin
        _zz_24_ <= (2'b00);
      end
      if(_zz_65_[24])begin
        _zz_25_ <= (2'b00);
      end
      if(_zz_65_[25])begin
        _zz_26_ <= (2'b00);
      end
      if(_zz_65_[26])begin
        _zz_27_ <= (2'b00);
      end
      if(_zz_65_[27])begin
        _zz_28_ <= (2'b00);
      end
      if(_zz_65_[28])begin
        _zz_29_ <= (2'b00);
      end
      if(_zz_65_[29])begin
        _zz_30_ <= (2'b00);
      end
      if(_zz_65_[30])begin
        _zz_31_ <= (2'b00);
      end
      if(_zz_65_[31])begin
        _zz_32_ <= (2'b00);
      end
      if(_zz_65_[32])begin
        _zz_33_ <= (2'b00);
      end
      if(_zz_65_[33])begin
        _zz_34_ <= (2'b00);
      end
      if(_zz_65_[34])begin
        _zz_35_ <= (2'b00);
      end
      if(_zz_65_[35])begin
        _zz_36_ <= (2'b00);
      end
      if(_zz_65_[36])begin
        _zz_37_ <= (2'b00);
      end
      if(_zz_65_[37])begin
        _zz_38_ <= (2'b00);
      end
      if(_zz_65_[38])begin
        _zz_39_ <= (2'b00);
      end
      if(_zz_65_[39])begin
        _zz_40_ <= (2'b00);
      end
      if(_zz_65_[40])begin
        _zz_41_ <= (2'b00);
      end
      if(_zz_65_[41])begin
        _zz_42_ <= (2'b00);
      end
      if(_zz_65_[42])begin
        _zz_43_ <= (2'b00);
      end
      if(_zz_65_[43])begin
        _zz_44_ <= (2'b00);
      end
      if(_zz_65_[44])begin
        _zz_45_ <= (2'b00);
      end
      if(_zz_65_[45])begin
        _zz_46_ <= (2'b00);
      end
      if(_zz_65_[46])begin
        _zz_47_ <= (2'b00);
      end
      if(_zz_65_[47])begin
        _zz_48_ <= (2'b00);
      end
      if(_zz_65_[48])begin
        _zz_49_ <= (2'b00);
      end
      if(_zz_65_[49])begin
        _zz_50_ <= (2'b00);
      end
      if(_zz_65_[50])begin
        _zz_51_ <= (2'b00);
      end
      if(_zz_65_[51])begin
        _zz_52_ <= (2'b00);
      end
      if(_zz_65_[52])begin
        _zz_53_ <= (2'b00);
      end
      if(_zz_65_[53])begin
        _zz_54_ <= (2'b00);
      end
      if(_zz_65_[54])begin
        _zz_55_ <= (2'b00);
      end
      if(_zz_65_[55])begin
        _zz_56_ <= (2'b00);
      end
      if(_zz_65_[56])begin
        _zz_57_ <= (2'b00);
      end
      if(_zz_65_[57])begin
        _zz_58_ <= (2'b00);
      end
      if(_zz_65_[58])begin
        _zz_59_ <= (2'b00);
      end
      if(_zz_65_[59])begin
        _zz_60_ <= (2'b00);
      end
      if(_zz_65_[60])begin
        _zz_61_ <= (2'b00);
      end
      if(_zz_65_[61])begin
        _zz_62_ <= (2'b00);
      end
      if(_zz_65_[62])begin
        _zz_63_ <= (2'b00);
      end
      if(_zz_65_[63])begin
        _zz_64_ <= (2'b00);
      end
    end
    if(wen_1)begin
      if(_zz_66_[0])begin
        _zz_1_ <= _zz_67_;
      end
      if(_zz_66_[1])begin
        _zz_2_ <= _zz_67_;
      end
      if(_zz_66_[2])begin
        _zz_3_ <= _zz_67_;
      end
      if(_zz_66_[3])begin
        _zz_4_ <= _zz_67_;
      end
      if(_zz_66_[4])begin
        _zz_5_ <= _zz_67_;
      end
      if(_zz_66_[5])begin
        _zz_6_ <= _zz_67_;
      end
      if(_zz_66_[6])begin
        _zz_7_ <= _zz_67_;
      end
      if(_zz_66_[7])begin
        _zz_8_ <= _zz_67_;
      end
      if(_zz_66_[8])begin
        _zz_9_ <= _zz_67_;
      end
      if(_zz_66_[9])begin
        _zz_10_ <= _zz_67_;
      end
      if(_zz_66_[10])begin
        _zz_11_ <= _zz_67_;
      end
      if(_zz_66_[11])begin
        _zz_12_ <= _zz_67_;
      end
      if(_zz_66_[12])begin
        _zz_13_ <= _zz_67_;
      end
      if(_zz_66_[13])begin
        _zz_14_ <= _zz_67_;
      end
      if(_zz_66_[14])begin
        _zz_15_ <= _zz_67_;
      end
      if(_zz_66_[15])begin
        _zz_16_ <= _zz_67_;
      end
      if(_zz_66_[16])begin
        _zz_17_ <= _zz_67_;
      end
      if(_zz_66_[17])begin
        _zz_18_ <= _zz_67_;
      end
      if(_zz_66_[18])begin
        _zz_19_ <= _zz_67_;
      end
      if(_zz_66_[19])begin
        _zz_20_ <= _zz_67_;
      end
      if(_zz_66_[20])begin
        _zz_21_ <= _zz_67_;
      end
      if(_zz_66_[21])begin
        _zz_22_ <= _zz_67_;
      end
      if(_zz_66_[22])begin
        _zz_23_ <= _zz_67_;
      end
      if(_zz_66_[23])begin
        _zz_24_ <= _zz_67_;
      end
      if(_zz_66_[24])begin
        _zz_25_ <= _zz_67_;
      end
      if(_zz_66_[25])begin
        _zz_26_ <= _zz_67_;
      end
      if(_zz_66_[26])begin
        _zz_27_ <= _zz_67_;
      end
      if(_zz_66_[27])begin
        _zz_28_ <= _zz_67_;
      end
      if(_zz_66_[28])begin
        _zz_29_ <= _zz_67_;
      end
      if(_zz_66_[29])begin
        _zz_30_ <= _zz_67_;
      end
      if(_zz_66_[30])begin
        _zz_31_ <= _zz_67_;
      end
      if(_zz_66_[31])begin
        _zz_32_ <= _zz_67_;
      end
      if(_zz_66_[32])begin
        _zz_33_ <= _zz_67_;
      end
      if(_zz_66_[33])begin
        _zz_34_ <= _zz_67_;
      end
      if(_zz_66_[34])begin
        _zz_35_ <= _zz_67_;
      end
      if(_zz_66_[35])begin
        _zz_36_ <= _zz_67_;
      end
      if(_zz_66_[36])begin
        _zz_37_ <= _zz_67_;
      end
      if(_zz_66_[37])begin
        _zz_38_ <= _zz_67_;
      end
      if(_zz_66_[38])begin
        _zz_39_ <= _zz_67_;
      end
      if(_zz_66_[39])begin
        _zz_40_ <= _zz_67_;
      end
      if(_zz_66_[40])begin
        _zz_41_ <= _zz_67_;
      end
      if(_zz_66_[41])begin
        _zz_42_ <= _zz_67_;
      end
      if(_zz_66_[42])begin
        _zz_43_ <= _zz_67_;
      end
      if(_zz_66_[43])begin
        _zz_44_ <= _zz_67_;
      end
      if(_zz_66_[44])begin
        _zz_45_ <= _zz_67_;
      end
      if(_zz_66_[45])begin
        _zz_46_ <= _zz_67_;
      end
      if(_zz_66_[46])begin
        _zz_47_ <= _zz_67_;
      end
      if(_zz_66_[47])begin
        _zz_48_ <= _zz_67_;
      end
      if(_zz_66_[48])begin
        _zz_49_ <= _zz_67_;
      end
      if(_zz_66_[49])begin
        _zz_50_ <= _zz_67_;
      end
      if(_zz_66_[50])begin
        _zz_51_ <= _zz_67_;
      end
      if(_zz_66_[51])begin
        _zz_52_ <= _zz_67_;
      end
      if(_zz_66_[52])begin
        _zz_53_ <= _zz_67_;
      end
      if(_zz_66_[53])begin
        _zz_54_ <= _zz_67_;
      end
      if(_zz_66_[54])begin
        _zz_55_ <= _zz_67_;
      end
      if(_zz_66_[55])begin
        _zz_56_ <= _zz_67_;
      end
      if(_zz_66_[56])begin
        _zz_57_ <= _zz_67_;
      end
      if(_zz_66_[57])begin
        _zz_58_ <= _zz_67_;
      end
      if(_zz_66_[58])begin
        _zz_59_ <= _zz_67_;
      end
      if(_zz_66_[59])begin
        _zz_60_ <= _zz_67_;
      end
      if(_zz_66_[60])begin
        _zz_61_ <= _zz_67_;
      end
      if(_zz_66_[61])begin
        _zz_62_ <= _zz_67_;
      end
      if(_zz_66_[62])begin
        _zz_63_ <= _zz_67_;
      end
      if(_zz_66_[63])begin
        _zz_64_ <= _zz_67_;
      end
    end
    if(wen_2)begin
      if(_zz_68_[0])begin
        _zz_1_ <= _zz_69_;
      end
      if(_zz_68_[1])begin
        _zz_2_ <= _zz_69_;
      end
      if(_zz_68_[2])begin
        _zz_3_ <= _zz_69_;
      end
      if(_zz_68_[3])begin
        _zz_4_ <= _zz_69_;
      end
      if(_zz_68_[4])begin
        _zz_5_ <= _zz_69_;
      end
      if(_zz_68_[5])begin
        _zz_6_ <= _zz_69_;
      end
      if(_zz_68_[6])begin
        _zz_7_ <= _zz_69_;
      end
      if(_zz_68_[7])begin
        _zz_8_ <= _zz_69_;
      end
      if(_zz_68_[8])begin
        _zz_9_ <= _zz_69_;
      end
      if(_zz_68_[9])begin
        _zz_10_ <= _zz_69_;
      end
      if(_zz_68_[10])begin
        _zz_11_ <= _zz_69_;
      end
      if(_zz_68_[11])begin
        _zz_12_ <= _zz_69_;
      end
      if(_zz_68_[12])begin
        _zz_13_ <= _zz_69_;
      end
      if(_zz_68_[13])begin
        _zz_14_ <= _zz_69_;
      end
      if(_zz_68_[14])begin
        _zz_15_ <= _zz_69_;
      end
      if(_zz_68_[15])begin
        _zz_16_ <= _zz_69_;
      end
      if(_zz_68_[16])begin
        _zz_17_ <= _zz_69_;
      end
      if(_zz_68_[17])begin
        _zz_18_ <= _zz_69_;
      end
      if(_zz_68_[18])begin
        _zz_19_ <= _zz_69_;
      end
      if(_zz_68_[19])begin
        _zz_20_ <= _zz_69_;
      end
      if(_zz_68_[20])begin
        _zz_21_ <= _zz_69_;
      end
      if(_zz_68_[21])begin
        _zz_22_ <= _zz_69_;
      end
      if(_zz_68_[22])begin
        _zz_23_ <= _zz_69_;
      end
      if(_zz_68_[23])begin
        _zz_24_ <= _zz_69_;
      end
      if(_zz_68_[24])begin
        _zz_25_ <= _zz_69_;
      end
      if(_zz_68_[25])begin
        _zz_26_ <= _zz_69_;
      end
      if(_zz_68_[26])begin
        _zz_27_ <= _zz_69_;
      end
      if(_zz_68_[27])begin
        _zz_28_ <= _zz_69_;
      end
      if(_zz_68_[28])begin
        _zz_29_ <= _zz_69_;
      end
      if(_zz_68_[29])begin
        _zz_30_ <= _zz_69_;
      end
      if(_zz_68_[30])begin
        _zz_31_ <= _zz_69_;
      end
      if(_zz_68_[31])begin
        _zz_32_ <= _zz_69_;
      end
      if(_zz_68_[32])begin
        _zz_33_ <= _zz_69_;
      end
      if(_zz_68_[33])begin
        _zz_34_ <= _zz_69_;
      end
      if(_zz_68_[34])begin
        _zz_35_ <= _zz_69_;
      end
      if(_zz_68_[35])begin
        _zz_36_ <= _zz_69_;
      end
      if(_zz_68_[36])begin
        _zz_37_ <= _zz_69_;
      end
      if(_zz_68_[37])begin
        _zz_38_ <= _zz_69_;
      end
      if(_zz_68_[38])begin
        _zz_39_ <= _zz_69_;
      end
      if(_zz_68_[39])begin
        _zz_40_ <= _zz_69_;
      end
      if(_zz_68_[40])begin
        _zz_41_ <= _zz_69_;
      end
      if(_zz_68_[41])begin
        _zz_42_ <= _zz_69_;
      end
      if(_zz_68_[42])begin
        _zz_43_ <= _zz_69_;
      end
      if(_zz_68_[43])begin
        _zz_44_ <= _zz_69_;
      end
      if(_zz_68_[44])begin
        _zz_45_ <= _zz_69_;
      end
      if(_zz_68_[45])begin
        _zz_46_ <= _zz_69_;
      end
      if(_zz_68_[46])begin
        _zz_47_ <= _zz_69_;
      end
      if(_zz_68_[47])begin
        _zz_48_ <= _zz_69_;
      end
      if(_zz_68_[48])begin
        _zz_49_ <= _zz_69_;
      end
      if(_zz_68_[49])begin
        _zz_50_ <= _zz_69_;
      end
      if(_zz_68_[50])begin
        _zz_51_ <= _zz_69_;
      end
      if(_zz_68_[51])begin
        _zz_52_ <= _zz_69_;
      end
      if(_zz_68_[52])begin
        _zz_53_ <= _zz_69_;
      end
      if(_zz_68_[53])begin
        _zz_54_ <= _zz_69_;
      end
      if(_zz_68_[54])begin
        _zz_55_ <= _zz_69_;
      end
      if(_zz_68_[55])begin
        _zz_56_ <= _zz_69_;
      end
      if(_zz_68_[56])begin
        _zz_57_ <= _zz_69_;
      end
      if(_zz_68_[57])begin
        _zz_58_ <= _zz_69_;
      end
      if(_zz_68_[58])begin
        _zz_59_ <= _zz_69_;
      end
      if(_zz_68_[59])begin
        _zz_60_ <= _zz_69_;
      end
      if(_zz_68_[60])begin
        _zz_61_ <= _zz_69_;
      end
      if(_zz_68_[61])begin
        _zz_62_ <= _zz_69_;
      end
      if(_zz_68_[62])begin
        _zz_63_ <= _zz_69_;
      end
      if(_zz_68_[63])begin
        _zz_64_ <= _zz_69_;
      end
    end
    if(wen_3)begin
      if(_zz_70_[0])begin
        _zz_1_ <= _zz_71_;
      end
      if(_zz_70_[1])begin
        _zz_2_ <= _zz_71_;
      end
      if(_zz_70_[2])begin
        _zz_3_ <= _zz_71_;
      end
      if(_zz_70_[3])begin
        _zz_4_ <= _zz_71_;
      end
      if(_zz_70_[4])begin
        _zz_5_ <= _zz_71_;
      end
      if(_zz_70_[5])begin
        _zz_6_ <= _zz_71_;
      end
      if(_zz_70_[6])begin
        _zz_7_ <= _zz_71_;
      end
      if(_zz_70_[7])begin
        _zz_8_ <= _zz_71_;
      end
      if(_zz_70_[8])begin
        _zz_9_ <= _zz_71_;
      end
      if(_zz_70_[9])begin
        _zz_10_ <= _zz_71_;
      end
      if(_zz_70_[10])begin
        _zz_11_ <= _zz_71_;
      end
      if(_zz_70_[11])begin
        _zz_12_ <= _zz_71_;
      end
      if(_zz_70_[12])begin
        _zz_13_ <= _zz_71_;
      end
      if(_zz_70_[13])begin
        _zz_14_ <= _zz_71_;
      end
      if(_zz_70_[14])begin
        _zz_15_ <= _zz_71_;
      end
      if(_zz_70_[15])begin
        _zz_16_ <= _zz_71_;
      end
      if(_zz_70_[16])begin
        _zz_17_ <= _zz_71_;
      end
      if(_zz_70_[17])begin
        _zz_18_ <= _zz_71_;
      end
      if(_zz_70_[18])begin
        _zz_19_ <= _zz_71_;
      end
      if(_zz_70_[19])begin
        _zz_20_ <= _zz_71_;
      end
      if(_zz_70_[20])begin
        _zz_21_ <= _zz_71_;
      end
      if(_zz_70_[21])begin
        _zz_22_ <= _zz_71_;
      end
      if(_zz_70_[22])begin
        _zz_23_ <= _zz_71_;
      end
      if(_zz_70_[23])begin
        _zz_24_ <= _zz_71_;
      end
      if(_zz_70_[24])begin
        _zz_25_ <= _zz_71_;
      end
      if(_zz_70_[25])begin
        _zz_26_ <= _zz_71_;
      end
      if(_zz_70_[26])begin
        _zz_27_ <= _zz_71_;
      end
      if(_zz_70_[27])begin
        _zz_28_ <= _zz_71_;
      end
      if(_zz_70_[28])begin
        _zz_29_ <= _zz_71_;
      end
      if(_zz_70_[29])begin
        _zz_30_ <= _zz_71_;
      end
      if(_zz_70_[30])begin
        _zz_31_ <= _zz_71_;
      end
      if(_zz_70_[31])begin
        _zz_32_ <= _zz_71_;
      end
      if(_zz_70_[32])begin
        _zz_33_ <= _zz_71_;
      end
      if(_zz_70_[33])begin
        _zz_34_ <= _zz_71_;
      end
      if(_zz_70_[34])begin
        _zz_35_ <= _zz_71_;
      end
      if(_zz_70_[35])begin
        _zz_36_ <= _zz_71_;
      end
      if(_zz_70_[36])begin
        _zz_37_ <= _zz_71_;
      end
      if(_zz_70_[37])begin
        _zz_38_ <= _zz_71_;
      end
      if(_zz_70_[38])begin
        _zz_39_ <= _zz_71_;
      end
      if(_zz_70_[39])begin
        _zz_40_ <= _zz_71_;
      end
      if(_zz_70_[40])begin
        _zz_41_ <= _zz_71_;
      end
      if(_zz_70_[41])begin
        _zz_42_ <= _zz_71_;
      end
      if(_zz_70_[42])begin
        _zz_43_ <= _zz_71_;
      end
      if(_zz_70_[43])begin
        _zz_44_ <= _zz_71_;
      end
      if(_zz_70_[44])begin
        _zz_45_ <= _zz_71_;
      end
      if(_zz_70_[45])begin
        _zz_46_ <= _zz_71_;
      end
      if(_zz_70_[46])begin
        _zz_47_ <= _zz_71_;
      end
      if(_zz_70_[47])begin
        _zz_48_ <= _zz_71_;
      end
      if(_zz_70_[48])begin
        _zz_49_ <= _zz_71_;
      end
      if(_zz_70_[49])begin
        _zz_50_ <= _zz_71_;
      end
      if(_zz_70_[50])begin
        _zz_51_ <= _zz_71_;
      end
      if(_zz_70_[51])begin
        _zz_52_ <= _zz_71_;
      end
      if(_zz_70_[52])begin
        _zz_53_ <= _zz_71_;
      end
      if(_zz_70_[53])begin
        _zz_54_ <= _zz_71_;
      end
      if(_zz_70_[54])begin
        _zz_55_ <= _zz_71_;
      end
      if(_zz_70_[55])begin
        _zz_56_ <= _zz_71_;
      end
      if(_zz_70_[56])begin
        _zz_57_ <= _zz_71_;
      end
      if(_zz_70_[57])begin
        _zz_58_ <= _zz_71_;
      end
      if(_zz_70_[58])begin
        _zz_59_ <= _zz_71_;
      end
      if(_zz_70_[59])begin
        _zz_60_ <= _zz_71_;
      end
      if(_zz_70_[60])begin
        _zz_61_ <= _zz_71_;
      end
      if(_zz_70_[61])begin
        _zz_62_ <= _zz_71_;
      end
      if(_zz_70_[62])begin
        _zz_63_ <= _zz_71_;
      end
      if(_zz_70_[63])begin
        _zz_64_ <= _zz_71_;
      end
    end
  end

endmodule
