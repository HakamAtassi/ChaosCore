`default_nettype none
`timescale 1ns/100ps


module sim;

    initial $display("Running ChaosCore sim");




endmodule;